/*              %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
                %                                                                            %
                %          IMPLEMENTAÇÃO DE UMA TABELA VERDADE COM 3 BITS DE ENTRADA         %
                %                                                                            %
                %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
=============================================================================================================================
Autor: Telmo Paes
Data: 24/07/2023
=============================================================================================================================
Descrição:



=============================================================================================================================
*/

module truth_table_case(
  a,
  b,
  c,
  s);

  // Declaração de entradas e saídas:

  input a;
  input b;
  input c;
  output f;

  // Declaração de wires (sinais):

  wire a;
  wire b;
  wire c;

  // Declaração de variáveis:
  
  reg s;

  // Inicia a rotina sequencial:
  
  always @(a or b or c)
  begin
    case({a,b,c})
      3'b000    :    s = 0;
      3'b001    :    s = 0;
      3'b010    :    s = 1;  
      3'b011    :    s = 1;
      3'b100    :    s = 0;
      3'b101    :    s = 0;
      3'b110    :    s = 1;
      3'b111    :    s = 0;
    endcase
  end
        
end module

  
